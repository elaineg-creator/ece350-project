module cpgenerate(g,p,a,b);

    input  [31:0] a,b;

    output [31:0] g,p;

    cla_slice s0(g[0],p[0],a[0],b[0]);

    cla_slice s1(g[1],p[1],a[1],b[1]);

    cla_slice s2(g[2],p[2],a[2],b[2]);

    cla_slice s3(g[3],p[3],a[3],b[3]);

    cla_slice s4(g[4],p[4],a[4],b[4]);

    cla_slice s5(g[5],p[5],a[5],b[5]);

    cla_slice s6(g[6],p[6],a[6],b[6]);

    cla_slice s7(g[7],p[7],a[7],b[7]);

    cla_slice s8(g[8],p[8],a[8],b[8]);

    cla_slice s9(g[9],p[9],a[9],b[9]);

    cla_slice s10(g[10],p[10],a[10],b[10]);

    cla_slice s11(g[11],p[11],a[11],b[11]);

    cla_slice s12(g[12],p[12],a[12],b[12]);

    cla_slice s13(g[13],p[13],a[13],b[13]);

    cla_slice s14(g[14],p[14],a[14],b[14]);

    cla_slice s15(g[15],p[15],a[15],b[15]);

    cla_slice s16(g[16],p[16],a[16],b[16]);

    cla_slice s17(g[17],p[17],a[17],b[17]);

    cla_slice s18(g[18],p[18],a[18],b[18]);

    cla_slice s19(g[19],p[19],a[19],b[19]);

    cla_slice s20(g[20],p[20],a[20],b[20]);

    cla_slice s21(g[21],p[21],a[21],b[21]);

    cla_slice s22(g[22],p[22],a[22],b[22]);

    cla_slice s23(g[23],p[23],a[23],b[23]);

    cla_slice s24(g[24],p[24],a[24],b[24]);

    cla_slice s25(g[25],p[25],a[25],b[25]);

    cla_slice s26(g[26],p[26],a[26],b[26]);

    cla_slice s27(g[27],p[27],a[27],b[27]);

    cla_slice s28(g[28],p[28],a[28],b[28]);

    cla_slice s29(g[29],p[29],a[29],b[29]);

    cla_slice s30(g[30],p[30],a[30],b[30]);

    cla_slice s31(g[31],p[31],a[31],b[31]);

 

endmodule