module bitwise_not(a, out);
    input [31:0] a;
    output [31:0] out;

    not NOT0(out[0], a[0]);
    not NOT1(out[1], a[1]);
    not NOT2(out[2], a[2]);
    not NOT3(out[3], a[3]);
    not NOT4(out[4], a[4]);
    not NOT5(out[5], a[5]);
    not NOT6(out[6], a[6]);
    not NOT7(out[7], a[7]);
    not NOT8(out[8], a[8]);
    not NOT9(out[9], a[9]);
    not NOT10(out[10], a[10]);
    not NOT11(out[11], a[11]);
    not NOT12(out[12], a[12]);
    not NOT13(out[13], a[13]);
    not NOT14(out[14], a[14]);
    not NOT15(out[15], a[15]);
    not NOT16(out[16], a[16]);
    not NOT17(out[17], a[17]);
    not NOT18(out[18], a[18]);
    not NOT19(out[19], a[19]);
    not NOT20(out[20], a[20]);
    not NOT21(out[21], a[21]);
    not NOT22(out[22], a[22]);
    not NOT23(out[23], a[23]);
    not NOT24(out[24], a[24]);
    not NOT25(out[25], a[25]);
    not NOT26(out[26], a[26]);
    not NOT27(out[27], a[27]);
    not NOT28(out[28], a[28]);
    not NOT29(out[29], a[29]);
    not NOT30(out[30], a[30]);
    not NOT31(out[31], a[31]);

    
endmodule