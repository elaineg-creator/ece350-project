module bitwise_and(a, b, out);
    input [31:0] a, b;
    output [31:0] out;

    and AND0(out[0], a[0], b[0]);
    and AND1(out[1], a[1], b[1]);
    and AND2(out[2], a[2], b[2]);
    and AND3(out[3], a[3], b[3]);
    and AND4(out[4], a[4], b[4]);
    and AND5(out[5], a[5], b[5]);
    and AND6(out[6], a[6], b[6]);
    and AND7(out[7], a[7], b[7]);
    and AND8(out[8], a[8], b[8]);
    and AND9(out[9], a[9], b[9]);
    and AND10(out[10], a[10], b[10]);
    and AND11(out[11], a[11], b[11]);
    and AND12(out[12], a[12], b[12]);
    and AND13(out[13], a[13], b[13]);
    and AND14(out[14], a[14], b[14]);
    and AND15(out[15], a[15], b[15]);
    and AND16(out[16], a[16], b[16]);
    and AND17(out[17], a[17], b[17]);
    and AND18(out[18], a[18], b[18]);
    and AND19(out[19], a[19], b[19]);
    and AND20(out[20], a[20], b[20]);
    and AND21(out[21], a[21], b[21]);
    and AND22(out[22], a[22], b[22]);
    and AND23(out[23], a[23], b[23]);
    and AND24(out[24], a[24], b[24]);
    and AND25(out[25], a[25], b[25]);
    and AND26(out[26], a[26], b[26]);
    and AND27(out[27], a[27], b[27]);
    and AND28(out[28], a[28], b[28]);
    and AND29(out[29], a[29], b[29]);
    and AND30(out[30], a[30], b[30]);
    and AND31(out[31], a[31], b[31]);

endmodule